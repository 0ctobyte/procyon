/* 
 * Copyright (c) 2019 Sekhar Bhattacharya
 *
 * SPDS-License-Identifier: MIT
 */

// Procyon constants

// ROB op types
`define PCYN_ROB_OP_WIDTH 2
`define PCYN_ROB_OP_INT   (`PCYN_ROB_OP_WIDTH'b00)
`define PCYN_ROB_OP_BR    (`PCYN_ROB_OP_WIDTH'b01)
`define PCYN_ROB_OP_LD    (`PCYN_ROB_OP_WIDTH'b10)
`define PCYN_ROB_OP_ST    (`PCYN_ROB_OP_WIDTH'b11)

// General operation types according to RV spec
`define PCYN_OPCODE_WIDTH  7
`define PCYN_OPCODE_OPIMM  (`PCYN_OPCODE_WIDTH'b0010011)
`define PCYN_OPCODE_LUI    (`PCYN_OPCODE_WIDTH'b0110111)
`define PCYN_OPCODE_AUIPC  (`PCYN_OPCODE_WIDTH'b0010111)
`define PCYN_OPCODE_OP     (`PCYN_OPCODE_WIDTH'b0110011)
`define PCYN_OPCODE_JAL    (`PCYN_OPCODE_WIDTH'b1101111)
`define PCYN_OPCODE_JALR   (`PCYN_OPCODE_WIDTH'b1100111)
`define PCYN_OPCODE_BRANCH (`PCYN_OPCODE_WIDTH'b1100011)
`define PCYN_OPCODE_LOAD   (`PCYN_OPCODE_WIDTH'b0000011)
`define PCYN_OPCODE_STORE  (`PCYN_OPCODE_WIDTH'b0100011)

// ALU operations
`define PCYN_ALU_FUNC_WIDTH  4
`define PCYN_ALU_SHAMT_WIDTH 5
`define PCYN_ALU_FUNC_ADD    (`PCYN_ALU_FUNC_WIDTH'b0000)
`define PCYN_ALU_FUNC_SUB    (`PCYN_ALU_FUNC_WIDTH'b0001)
`define PCYN_ALU_FUNC_AND    (`PCYN_ALU_FUNC_WIDTH'b0010)
`define PCYN_ALU_FUNC_OR     (`PCYN_ALU_FUNC_WIDTH'b0011)
`define PCYN_ALU_FUNC_XOR    (`PCYN_ALU_FUNC_WIDTH'b0100)
`define PCYN_ALU_FUNC_SLL    (`PCYN_ALU_FUNC_WIDTH'b0101)
`define PCYN_ALU_FUNC_SRL    (`PCYN_ALU_FUNC_WIDTH'b0110)
`define PCYN_ALU_FUNC_SRA    (`PCYN_ALU_FUNC_WIDTH'b0111)
`define PCYN_ALU_FUNC_EQ     (`PCYN_ALU_FUNC_WIDTH'b1000)
`define PCYN_ALU_FUNC_NE     (`PCYN_ALU_FUNC_WIDTH'b1001)
`define PCYN_ALU_FUNC_LT     (`PCYN_ALU_FUNC_WIDTH'b1010)
`define PCYN_ALU_FUNC_LTU    (`PCYN_ALU_FUNC_WIDTH'b1011)
`define PCYN_ALU_FUNC_GE     (`PCYN_ALU_FUNC_WIDTH'b1100)
`define PCYN_ALU_FUNC_GEU    (`PCYN_ALU_FUNC_WIDTH'b1101)

// LSU operations
`define PCYN_LSU_FUNC_WIDTH 4
`define PCYN_LSU_FUNC_LB    (`PCYN_LSU_FUNC_WIDTH'b0000)
`define PCYN_LSU_FUNC_LH    (`PCYN_LSU_FUNC_WIDTH'b0001)
`define PCYN_LSU_FUNC_LW    (`PCYN_LSU_FUNC_WIDTH'b0010)
`define PCYN_LSU_FUNC_LBU   (`PCYN_LSU_FUNC_WIDTH'b0011)
`define PCYN_LSU_FUNC_LHU   (`PCYN_LSU_FUNC_WIDTH'b0100)
`define PCYN_LSU_FUNC_SB    (`PCYN_LSU_FUNC_WIDTH'b0101)
`define PCYN_LSU_FUNC_SH    (`PCYN_LSU_FUNC_WIDTH'b0110)
`define PCYN_LSU_FUNC_SW    (`PCYN_LSU_FUNC_WIDTH'b0111)
`define PCYN_LSU_FUNC_FILL  (`PCYN_LSU_FUNC_WIDTH'b1000)

// BIU operations
`define PCYN_BIU_FUNC_WIDTH 2
`define PCYN_BIU_FUNC_READ  (`PCYN_BIU_FUNC_WIDTH'b00)
`define PCYN_BIU_FUNC_WRITE (`PCYN_BIU_FUNC_WIDTH'b01)
`define PCYN_BIU_FUNC_RMW   (`PCYN_BIU_FUNC_WIDTH'b10)

// BIU burst lengths
`define PCYN_BIU_LEN_WIDTH    3
`define PCYN_BIU_LEN_1B       (`PCYN_BIU_LEN_WIDTH'b000)
`define PCYN_BIU_LEN_2B       (`PCYN_BIU_LEN_WIDTH'b001)
`define PCYN_BIU_LEN_4B       (`PCYN_BIU_LEN_WIDTH'b010)
`define PCYN_BIU_LEN_8B       (`PCYN_BIU_LEN_WIDTH'b011)
`define PCYN_BIU_LEN_16B      (`PCYN_BIU_LEN_WIDTH'b100)
`define PCYN_BIU_LEN_32B      (`PCYN_BIU_LEN_WIDTH'b101)
`define PCYN_BIU_LEN_64B      (`PCYN_BIU_LEN_WIDTH'b110)
`define PCYN_BIU_LEN_128B     (`PCYN_BIU_LEN_WIDTH'b111)
`define PCYN_BIU_LEN_MAX      (`PCYN_BIU_LEN_128B)
`define PCYN_BIU_LEN_MAX_SIZE 128

// Wishbone bus Cycle Type Identifiers
`define WB_CTI_WIDTH        3
`define WB_CTI_CLASSIC      (`WB_CTI_WIDTH'b000)
`define WB_CTI_CONSTANT     (`WB_CTI_WIDTH'b001)
`define WB_CTI_INCREMENTING (`WB_CTI_WIDTH'b010)
`define WB_CTI_END_OF_BURST (`WB_CTI_WIDTH'b111)

// Wishbone bus Burst Type Extensions
`define WB_BTE_WIDTH 2
`define WB_BTE_LINEAR (`WB_BTE_WIDTH'b00)
`define WB_BTE_4BEAT  (`WB_BTE_WIDTH'b01)
`define WB_BTE_8BEAT  (`WB_BTE_WIDTH'b10)
`define WB_BTE_16BEAT (`WB_BTE_WIDTH'b11)
