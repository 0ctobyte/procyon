// Procyon constants

// ROB op types
`define PCYN_ROB_OP_WIDTH 2
`define PCYN_ROB_OP_INT   (`PCYN_ROB_OP_WIDTH'b00)
`define PCYN_ROB_OP_BR    (`PCYN_ROB_OP_WIDTH'b01)
`define PCYN_ROB_OP_LD    (`PCYN_ROB_OP_WIDTH'b10)
`define PCYN_ROB_OP_ST    (`PCYN_ROB_OP_WIDTH'b11)

// General operation types according to RV spec
`define PCYN_OPCODE_WIDTH  7
`define PCYN_OPCODE_OPIMM  (`PCYN_OPCODE_WIDTH'b0010011)
`define PCYN_OPCODE_LUI    (`PCYN_OPCODE_WIDTH'b0110111)
`define PCYN_OPCODE_AUIPC  (`PCYN_OPCODE_WIDTH'b0010111)
`define PCYN_OPCODE_OP     (`PCYN_OPCODE_WIDTH'b0110011)
`define PCYN_OPCODE_JAL    (`PCYN_OPCODE_WIDTH'b1101111)
`define PCYN_OPCODE_JALR   (`PCYN_OPCODE_WIDTH'b1100111)
`define PCYN_OPCODE_BRANCH (`PCYN_OPCODE_WIDTH'b1100011)
`define PCYN_OPCODE_LOAD   (`PCYN_OPCODE_WIDTH'b0000011)
`define PCYN_OPCODE_STORE  (`PCYN_OPCODE_WIDTH'b0100011)

// ALU operations
`define PCYN_ALU_FUNC_WIDTH  4
`define PCYN_ALU_SHAMT_WIDTH 5
`define PCYN_ALU_FUNC_ADD    (`PCYN_ALU_FUNC_WIDTH'b0000)
`define PCYN_ALU_FUNC_SUB    (`PCYN_ALU_FUNC_WIDTH'b0001)
`define PCYN_ALU_FUNC_AND    (`PCYN_ALU_FUNC_WIDTH'b0010)
`define PCYN_ALU_FUNC_OR     (`PCYN_ALU_FUNC_WIDTH'b0011)
`define PCYN_ALU_FUNC_XOR    (`PCYN_ALU_FUNC_WIDTH'b0100)
`define PCYN_ALU_FUNC_SLL    (`PCYN_ALU_FUNC_WIDTH'b0101)
`define PCYN_ALU_FUNC_SRL    (`PCYN_ALU_FUNC_WIDTH'b0110)
`define PCYN_ALU_FUNC_SRA    (`PCYN_ALU_FUNC_WIDTH'b0111)
`define PCYN_ALU_FUNC_EQ     (`PCYN_ALU_FUNC_WIDTH'b1000)
`define PCYN_ALU_FUNC_NE     (`PCYN_ALU_FUNC_WIDTH'b1001)
`define PCYN_ALU_FUNC_LT     (`PCYN_ALU_FUNC_WIDTH'b1010)
`define PCYN_ALU_FUNC_LTU    (`PCYN_ALU_FUNC_WIDTH'b1011)
`define PCYN_ALU_FUNC_GE     (`PCYN_ALU_FUNC_WIDTH'b1100)
`define PCYN_ALU_FUNC_GEU    (`PCYN_ALU_FUNC_WIDTH'b1101)

// LSU operations
`define PCYN_LSU_FUNC_WIDTH 4
`define PCYN_LSU_FUNC_LB    (`PCYN_LSU_FUNC_WIDTH'b0000)
`define PCYN_LSU_FUNC_LH    (`PCYN_LSU_FUNC_WIDTH'b0001)
`define PCYN_LSU_FUNC_LW    (`PCYN_LSU_FUNC_WIDTH'b0010)
`define PCYN_LSU_FUNC_LBU   (`PCYN_LSU_FUNC_WIDTH'b0011)
`define PCYN_LSU_FUNC_LHU   (`PCYN_LSU_FUNC_WIDTH'b0100)
`define PCYN_LSU_FUNC_SB    (`PCYN_LSU_FUNC_WIDTH'b0101)
`define PCYN_LSU_FUNC_SH    (`PCYN_LSU_FUNC_WIDTH'b0110)
`define PCYN_LSU_FUNC_SW    (`PCYN_LSU_FUNC_WIDTH'b0111)
`define PCYN_LSU_FUNC_FILL  (`PCYN_LSU_FUNC_WIDTH'b1000)
